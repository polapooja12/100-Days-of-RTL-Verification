interface sub_inf;
    logic a;
    logic b;
    logic bin;
    bit diff;
    bit bout;
endinterface
