interface decoder_inf; // Interface for the decoder
    logic a; // Input a
    logic b; // Input b
    logic y0; // Output y0
    logic y1; // Output y1
    logic y2; // Output y2
    logic y3; // Output y3
endinterface
