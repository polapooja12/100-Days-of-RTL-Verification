interface clock_divider_inf;
    logic clk;  // Clock signal
    logic f2;   // Divided frequency signals
    logic f4;
    logic f8;
    logic f16;
    logic f32;
    logic f64;
endinterface
