interface sync_counter_inf;
    logic clk; 
    logic [3:0] q;      // Output from the synchronous counter
    logic [3:0] qbar;   // Inverted output from the synchronous counter
endinterface
