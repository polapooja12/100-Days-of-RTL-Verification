// sipo_interface.sv
interface sipo_inf;
    logic clk; 
    logic d; 
    logic [3:0] q; // Output from the SIPO register
endinterface
