interface rca_interface;
    logic [3:0] a, b;
    logic cin;
    logic [3:0] sum;
    logic carryout;
endinterface
