module comp(a,b,x,y,z);
 input wire a,b;
 output reg,y,2;
 assign x=-(a^b);//equal
 assign y=(-a&b);//lesser
  assign z= (a&~b);//greater
endmodule


