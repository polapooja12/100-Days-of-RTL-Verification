interface add_inf;
logic a;
logic b;
logic cin;
bit sum;
bit carry;
endinterface
