interface jk_ff_if;
    logic clk;    // Clock signal
    logic reset;  // Asynchronous reset signal
    logic j;      // J input
    logic k;      // K input
    logic q;      // Q output
    logic qn;     // Complementary Q output
endinterface
