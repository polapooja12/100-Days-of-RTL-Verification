interface BCDto7Segment_inf;
  logic [3:0] bcd;  // 4-bit BCD input
  logic [6:0] seg;  // 7-segment output (a-g)
endinterface
