interface full_inf; // Interface for the MUX
    logic a, b, c, d;   // 4 data inputs
    logic s1, s2;       // 2-bit select input
    logic y;            // Output
endinterface
