interface priority_encoder_if;
  logic a;   // Input a
  logic b;   // Input b
  logic c;   // Input c
  logic d;   // Input d
  logic y1;  // Output y1
  logic y2;  // Output y2
endinterface
