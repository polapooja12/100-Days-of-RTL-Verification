interface logicgates_inf;
  logic a;
  logic b;
  logic y1, y2, y3, y4, y5, y6;
endinterface
